`default_nettype none

module clk_wiz_0
  (
   output wire clk_out1,
   input  wire reset,
   output wire locked,
   input  wire clk_in1
   );

endmodule // clk_wiz_0

`default_nettype wire

